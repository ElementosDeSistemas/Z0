library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Mux4Way is
	port ( 
			a:   in  STD_LOGIC;
			b:   in  STD_LOGIC;
			c:   in  STD_LOGIC;
			d:   in  STD_LOGIC;
			sel: in  STD_LOGIC_VECTOR(1 downto 0);
			q:   out STD_LOGIC);
end entity;
	
	architecture Run of Mux4Way is
		begin
		with (sel) select
      q <= a when '00',
		q <= b when '01',
		q <= c when '10',
		q <= d when '11'
	end architecture;